`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:04:43 01/08/2017 
// Design Name: 
// Module Name:    HAHA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module HAHA(clk,row,col,haha
    );

input clk;
reg flag;
input [10:0]row,col;
output reg [2:0] haha;

wire [10:0]sr;
wire [299:0] r_1, r_2,r_3,r_4,r_5,r_6,r_7,r_8,r_9,r_10,r_11,r_12,r_13,r_14,r_15,r_16,r_17,r_18,r_19,r_20;
wire [299:0] r_21,r_22,r_23,r_24,r_25,r_26,r_27,r_28,r_29,r_30,r_31,r_32,r_33,r_34,r_35,r_36,r_37,r_38,r_39,r_40;
wire [299:0] r_41,r_42,r_43,r_44,r_45,r_46,r_47,r_48,r_49,r_50,r_51,r_52,r_53,r_54,r_55,r_56,r_57,r_58,r_59,r_60;
wire [299:0] r_61,r_62,r_63,r_64,r_65,r_66,r_67,r_68,r_69,r_70,r_71,r_72,r_73,r_74,r_75,r_76,r_77,r_78,r_79,r_80;
wire [299:0] r_81,r_82,r_83,r_84,r_85,r_86,r_87,r_88,r_89,r_90,r_91,r_92,r_93,r_94,r_95,r_96,r_97,r_98,r_99,r_100;
wire [299:0] r_101,r_102,r_103,r_104,r_105,r_106,r_107,r_108,r_109,r_110,r_111,r_112,r_113,r_114,r_115,r_116,r_117,r_118,r_119,r_120;
wire [299:0] r_121,r_122,r_123,r_124,r_125,r_126,r_127,r_128,r_129,r_130,r_131,r_132,r_133,r_134,r_135,r_136,r_137,r_138,r_139,r_140;
wire [299:0] r_141,r_142,r_143,r_144;

assign sr = row-50;

assign r_1   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_2   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_3   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_4   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_5   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000111111111110000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_6   = 200'b00000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000111111111110000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_7   = 200'b00000000000000000000000000000000000000000000000000000000000000000000111111111100000000000001111111111111111110000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_8   = 200'b00000000000000000000000000000000000000000000000000000000000000000000111111111100000000000001111111111111111110000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_9   = 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000000000000000111111000000000011111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000 ;
assign r_10  = 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000000000000000111111000000000011111100000000000000000111111100000000000000000000000000000000000000000000000000000000000000000 ;
assign r_11  = 200'b00000000000000000000000000000000000000000000000000000000000000111111100001111111110000001111000000000000000011110000000000000000000111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_12  = 200'b00000000000000000000000000000000000000000000000000000000000000111111100001111111110000001111000000000000000011110000000000000000000111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_13  = 200'b00000000000000000000000000000000000000000000000000000000010111111100011111111111111111011111111100000000000001111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000 ;
assign r_14  = 200'b00000000000000000000000000000000000000000000000000000000010111111100011111111111111111011111111100000000000001111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000 ;
assign r_15  = 200'b00000000000000000000000000000000000000000000000000000000111111100001111110000000111111111111111110000000000000111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000 ;
assign r_16  = 200'b00000000000000000000000000000000000000000000000000000000111111100001111110000000111111111111111110000000000000111100000000000000000000111111110000000000000000000000000000000000000000000000000000000000 ;
assign r_17  = 200'b00000000000000000000000000000000000000000000000000000011111110000011110000000000111111111111111110000000000000011111111100000000000000000011110000000000000000000000000000000000000000000000000000000000 ;
assign r_18  = 200'b00000000000000000000000000000000000000000000000000000011111110000011110000000000111111111111111110000000000000011111111100000000000000000011110000000000000000000000000000000000000000000000000000000000 ;
assign r_19  = 200'b00000000000000000000000000000000000000000000000000001111110000000111000000000000111111111111111100000000000000011111111111111111111111110001111100000000000000000000000000000000000000000000000000000000 ;
assign r_20  = 200'b00000000000000000000000000000000000000000000000000001111110000000111000000000000111111111111111100000000000000011111111111111111111111110001111100000000000000000000000000000000000000000000000000000000 ;
assign r_21  = 200'b00000000000000000000000000000000000000000000000000111111000000001110000000000000111111011110110000000000000000111100000011111111111111111110111110000000000000000000000000000000000000000000000000000000 ;
assign r_22  = 200'b00000000000000000000000000000000000000000000000000111111000000001110000000000000111111011110110000000000000000111100000011111111111111111110111110000000000000000000000000000000000000000000000000000000 ;
assign r_23  = 200'b00000000000000000000000000000000000000000000000001111100000000001110000000000000011111101110000000000000000000111000000001111110000000111111011111000000000000000000000000000000000000000000000000000000 ;
assign r_24  = 200'b00000000000000000000000000000000000000000000000001111100000000001110000000000000011111101110000000000000000000111000000001111110000000111111011111000000000000000000000000000000000000000000000000000000 ;
assign r_25  = 200'b00000000000000000000000000000000000000000000000111110000000000011100000000000000000000011111100000000000000011110011111000000000000000000111100111100000000000000000000000000000000000000000000000000000 ;
assign r_26  = 200'b00000000000000000000000000000000000000000000000111110000000000011100000000000000000000011111100000000000000011110011111000000000000000000111100111100000000000000000000000000000000000000000000000000000 ;
assign r_27  = 200'b00000000000000000000000000000000000000000000001111100000000000011100000000000000000000011111111110000000111111111111111000000000000000000011110011110000000000000000000000000000000000000000000000000000 ;
assign r_28  = 200'b00000000000000000000000000000000000000000000001111100000000000011100000000000000000000011111111110000000111111111111111000000000000000000011110011110000000000000000000000000000000000000000000000000000 ;
assign r_29  = 200'b00000000000000000000000000000000000000000000111110000000000000001110000000000000000001111111111111111111111111111110000000011000000000000001110001110000000000000000000000000000000000000000000000000000 ;
assign r_30  = 200'b00000000000000000000000000000000000000000000111110000000000000001110000000000000000001111111111111111111111111111110000000011000000000000001110001110000000000000000000000000000000000000000000000000000 ;
assign r_31  = 200'b00000000000000000000000000000000000000000000111100000000000011111111100000000000000011110011000011111111111111100000011111111100000000000001110001111000000000000000000000000000000000000000000000000000 ;
assign r_32  = 200'b00000000000000000000000000000000000000000000111100000000000011111111100000000000000011110011000011111111111111100000011111111100000000000001110001111000000000000000000000000000000000000000000000000000 ;
assign r_33  = 200'b00000000000000000000000000000000000000000001111000000000001111111111111000000000001111101000000011100111111100011111111111110000000000000011110000111100000000000000000000000000000000000000000000000000 ;
assign r_34  = 200'b00000000000000000000000000000000000000000001111000000000001111111111111000000000001111101000000011100111111100011111111111110000000000000011110000111100000000000000000000000000000000000000000000000000 ;
assign r_35  = 200'b00000000000000000000000000000000000000000011110000000000111111000001111111111111111111100000000111100001111111111111110000000100000000000011110000011110000000000000000000000000000000000000000000000000 ;
assign r_36  = 200'b00000000000000000000000000000000000000000011110000000000111111000001111111111111111111100000000111100001111111111111110000000100000000000011110000011110000000000000000000000000000000000000000000000000 ;
assign r_37  = 200'b00000000000000000000000000000000000000000111100000011111111100000011011111111111111111111111111111000000111111110001111111111110000000001111111100011110000000000000000000000000000000000000000000000000 ;
assign r_38  = 200'b00000000000000000000000000000000000000000111100000011111111100000011011111111111111111111111111111000000111111110001111111111110000000001111111100011110000000000000000000000000000000000000000000000000 ;
assign r_39  = 200'b00000000000000000000000000000000000000001111000001111111111111000011111111111111111110111111111100000000100111111111111111111100000000111110011110001110000000000000000000000000000000000000000000000000 ;
assign r_40  = 200'b00000000000000000000000000000000000000001111000001111111111111000011111111111111111110111111111100000000100111111111111111111100000000111110011110001110000000000000000000000000000000000000000000000000 ;
assign r_41  = 200'b00000000000000000000000000000000000000001110000111111010011110000001111111111111111100000011111000000000001111111111100000000000011111111100001110001110000000000000000000000000000000000000000000000000 ;
assign r_42  = 200'b00000000000000000000000000000000000000001110000111111010011110000001111111111111111100000011111000000000001111111111100000000000011111111100001110001110000000000000000000000000000000000000000000000000 ;
assign r_43  = 200'b00000000000000000000000000000000000000001110001111000000000000000000001111111111111111000000111100000000000100000000111111111111111111111000001111001110000000000000000000000000000000000000000000000000 ;
assign r_44  = 200'b00000000000000000000000000000000000000001110001111000000000000000000001111111111111111000000111100000000000100000000111111111111111111111000001111001110000000000000000000000000000000000000000000000000 ;
assign r_45  = 200'b00000000000000000000000000000000000000011110001110000000000000000111111111111111111111000000011100000000111111111111111111111111110000111000000011101111000000000000000000000000000000000000000000000000 ;
assign r_46  = 200'b00000000000000000000000000000000000000011110001110000000000000000111111111111111111111000000011100000000111111111111111111111111110000111000000011101111000000000000000000000000000000000000000000000000 ;
assign r_47  = 200'b00000000000000000000000000000000000000011100011100000000000000000011111110000011111111100000001111111111111111111111111000000000000000111000000011100111011111111110000000000000000000000000000000000000 ;
assign r_48  = 200'b00000000000000000000000000000000000000011100011100000000000000000011111110000011111111100000001111111111111111111111111000000000000000111000000011100111011111111110000000000000000000000000000000000000 ;
assign r_49  = 200'b00000000000000000000000000000000000000111100011100000000000000000000000111111111111111000111111111111111100000000000000000000000000000111000000001111111111111111111110000000000000000000000000000000000 ;
assign r_50  = 200'b00000000000000000000000000000000000000111100011100000000000000000000000111111111111111000111111111111111100000000000000000000000000000111000000001111111111111111111110000000000000000000000000000000000 ;
assign r_51  = 200'b00000000000000000000000000000000000000111100011100000000000000000011111111111111000011111111111110000000000000000000000000000000000000111000000001110111111000000011111000000000000000000000000000000000 ;
assign r_52  = 200'b00000000000000000000000000000000000000111100011100000000000000000011111111111111000011111111111110000000000000000000000000000000000000111000000001110111111000000011111000000000000000000000000000000000 ;
assign r_53  = 200'b00000000000000000000000000000000000000111000011110000000000000000011111111000001111111111100000000000000000000000000000000000000000000111000000001110111000000000000111110000000000000000000000000000000 ;
assign r_54  = 200'b00000000000000000000000000000000000000111000011110000000000000000011111111000001111111111100000000000000000000000000000000000000000000111000000001110111000000000000111110000000000000000000000000000000 ;
assign r_55  = 200'b00000000000000000000000000000000000000111100001111100000000000000000000000111111111110000000000000000000000000000000000000000000000000111000000001110111000000000000001110000000000000000000000000000000 ;
assign r_56  = 200'b00000000000000000000000000000000000000111100001111100000000000000000000000111111111110000000000000000000000000000000000000000000000000111000000001110111000000000000001110000000000000000000000000000000 ;
assign r_57  = 200'b00000000000000000000000000000000000000111100000111110000000000000000001111111111000000000000000000000000000000000000000000000000000001110000000001110111000000000000001111000111111111110000000000000000 ;
assign r_58  = 200'b00000000000000000000000000000000000000111100000111110000000000000000001111111111000000000000000000000000000000000000000000000000000001110000000001110111000000000000001111000111111111110000000000000000 ;
assign r_59  = 200'b00000000000000000000000000000000000000011100000011111111101001111111111111110000000000000000000000000000000000000000000000000000000001110000000001110111000000000000000111111111111111111111110000000000 ;
assign r_60  = 200'b00000000000000000000000000000000000000011100000011111111101001111111111111110000000000000000000000000000000000000000000000000000000001110000000001110111000000000000000111111111111111111111110000000000 ;
assign r_61  = 200'b00000000000000000000000000000000000000011100000111011111111111111111111000000000000000000000000000000000000000000000000000000000000011110000000001111111000000000000000111111110000000111111111110000000 ;
assign r_62  = 200'b00000000000000000000000000000000000000011100000111011111111111111111111000000000000000000000000000000000000000000000000000000000000011110000000001111111000000000000000111111110000000111111111110000000 ;
assign r_63  = 200'b00000000000000000000000000000000000000001110000111000000111111000000000000000000000000000000000000000000000000000000000000000000000011100000000001111110000000000000000111000000000000000000111111101000 ;
assign r_64  = 200'b00000000000000000000000000000000000000001110000111000000111111000000000000000000000000000000000000000000000000000000000000000000000011100000000001111110000000000000000111000000000000000000111111101000 ;
assign r_65  = 200'b00000000000000000000000000000000000000001110000111000000001111000000000000000000000000000000000000000000000000000000000000000000000011100000000001111110000000000000001111000000000000000000000111111000 ;
assign r_66  = 200'b00000000000000000000000000000000000000001110000111000000001111000000000000000000000000000000000000000000000000000000000000000000000011100000000001111110000000000000001111000000000000000000000111111000 ;
assign r_67  = 200'b00000000000000000000000000000000000000001111000111000000000111100000000000000000000000000000000000000000000000000000000000000000000111100000000001111100000000000000011110000011111111111111100000111110 ;
assign r_68  = 200'b00000000000000000000000000000000000000001111000111000000000111100000000000000000000000000000000000000000000000000000000000000000000111100000000001111100000000000000011110000011111111111111100000111110 ;
assign r_69  = 200'b00000000000000000000000000000000000000000111100111000000000011110000000000000000000000000000000000000000000000000000000000000000000111000000000011111100000000000000111111111111111111111111111111111111 ;
assign r_70  = 200'b00000000000000000000000000000000000000000111100111000000000011110000000000000000000000000000000000000000000000000000000000000000000111000000000011111100000000000000111111111111111111111111111111111111 ;
assign r_71  = 200'b00000000000000000000000000000000000000000011110111100000000001111000000000000000000000000000000000000000000000000011111111110000011110000000000011111000000000000001111111111111111000001111111111111111 ;
assign r_72  = 200'b00000000000000000000000000000000000000000011110111100000000001111000000000000000000000000000000000000000000000000011111111110000011110000000000011111000000000000001111111111111111000001111111111111111 ;
assign r_73  = 200'b00000000000000000000000000000000000000000001111011100000000000111100000000000000000000000000000000000000000000111111111111111111011100000000000111111100000000001111111001111000000000000000000000000000 ;
assign r_74  = 200'b00000000000000000000000000000000000000000001111011100000000000111100000000000000000000000000000000000000000000111111111111111111011100000000000111111100000000001111111001111000000000000000000000000000 ;
assign r_75  = 200'b00000000000000000000000000000000000011111111111101110000000000011111000000000000000000000000000000000000000111111110000000011111111100000000001111111111111111111111000001110000000000000000000000000000 ;
assign r_76  = 200'b00000000000000000000000000000000000011111111111101110000000000011111000000000000000000000000000000000000000111111110000000011111111100000000001111111111111111111111000001110000000000000000000000000000 ;
assign r_77  = 200'b00000000000000000000000000000000111111111111111111110000000000001111100000000000000000000111111111111111111111100000000000000011111000000000011111011111111111111100000011100000000000000000000000000000 ;
assign r_78  = 200'b00000000000000000000000000000000111111111111111111110000000000001111100000000000000000000111111111111111111111100000000000000011111000000000011111011111111111111100000011100000000000000000000000000000 ;
assign r_79  = 200'b00000000000000000000000000000011111111100111111111111100000000000011111000000000000000111111111111111111111000000000000000000011110000000000111110000001111110000000000111100000000000000000000000000000 ;
assign r_80  = 200'b00000000000000000000000000000011111111100111111111111100000000000011111000000000000000111111111111111111111000000000000000000011110000000000111110000001111110000000000111100000000000000000000000000000 ;
assign r_81  = 200'b00000000000000000000000000000111110000000000000111111100000000000001111110000000000011111100000000000000000000000000000000000111100000000011111100000001111000000000001111000000000000000000000000000000 ;
assign r_82  = 200'b00000000000000000000000000000111110000000000000111111100000000000001111110000000000011111100000000000000000000000000000000000111100000000011111100000001111000000000001111000000000000000000000000000000 ;
assign r_83  = 200'b00000000000000000000000000001111000000000000000011111110000000000000111111100000000111110000000000000000000000000000000000011110000000001111111000001111110000000000011110000000000000000000000000000000 ;
assign r_84  = 200'b00000000000000000000000000001111000000000000000011111110000000000000111111100000000111110000000000000000000000000000000000011110000000001111111000001111110000000000011110000000000000000000000000000000 ;
assign r_85  = 200'b00000000000000000000000000011110000000000000000001111111000000000000000111111000000111000000000000000000000000000000000001111100000000111111110000001111000000000000111100000000000000000000000000000000 ;
assign r_86  = 200'b00000000000000000000000000011110000000000000000001111111000000000000000111111000000111000000000000000000000000000000000001111100000000111111110000001111000000000000111100000000000000000000000000000000 ;
assign r_87  = 200'b00000000000000000000000000011100000000000000000000011111110000000000000000111111001110000000000000000000000000000000001111110000000011111111100000111110000000000001111000000000000000000000000000000000 ;
assign r_88  = 200'b00000000000000000000000000011100000000000000000000011111110000000000000000111111001110000000000000000000000000000000001111110000000011111111100000111110000000000001111000000000000000000000000000000000 ;
assign r_89  = 200'b00000000000000000000000000011100000000000000000000001111111000000000000000001111111100000000000000000000000000000001111111000000011111111111100011111100000000000011110000000000000000000000000000000000 ;
assign r_90  = 200'b00000000000000000000000000011100000000000000000000001111111000000000000000001111111100000000000000000000000000000001111111000000011111111111100011111100000000000011110000000000000000000000000000000000 ;
assign r_91  = 200'b00000000000000000000000000011100000000000000000000000001111110000000000000000001111111110000000000000000000000111111111000000001111111111111100111110000000000001111100000000000000000000000000000000000 ;
assign r_92  = 200'b00000000000000000000000000011100000000000000000000000001111110000000000000000001111111110000000000000000000000111111111000000001111111111111100111110000000000001111100000000000000000000000000000000000 ;
assign r_93  = 200'b00000000000000000000000000011110000000000000000000000001111111100000000000000000000111111111111111111111111111111110000000011111111111111111111111000000000001111110000000000000000000000000000000000000 ;
assign r_94  = 200'b00000000000000000000000000011110000000000000000000000001111111100000000000000000000111111111111111111111111111111110000000011111111111111111111111000000000001111110000000000000000000000000000000000000 ;
assign r_95  = 200'b00000000000000000000000000001110000000000000000000000001111111111100000000000000000000001111111111111111111111100000000111111111111111111111111100000000011111111000000000000000000000000000000000000000 ;
assign r_96  = 200'b00000000000000000000000000001110000000000000000000000001111111111100000000000000000000001111111111111111111111100000000111111111111111111111111100000000011111111000000000000000000000000000000000000000 ;
assign r_97  = 200'b00000000000000000000000000001111000000000000000000000011110001111111110000000000000000000000000000000000000000000011111111111011111111111111111111111111111111000000000000000000000000000000000000000000 ;
assign r_98  = 200'b00000000000000000000000000001111000000000000000000000011110001111111110000000000000000000000000000000000000000000011111111111011111111111111111111111111111111000000000000000000000000000000000000000000 ;
assign r_99  = 200'b00000000000000000000000000000111100000000000000000001111100000001111111111100000000000000000000000000000000011111111111110011111111111111000010111111111110000000000000000000000000000000000000000000000 ;
assign r_100 = 200'b00000000000000000000000000000111100000000000000000001111100000001111111111100000000000000000000000000000000011111111111110011111111111111000010111111111110000000000000000000000000000000000000000000000 ;
assign r_101 = 200'b00000000000000000000000111111111111100000000000000111111000000000011111111111111111110000000000001111111111111111111100111111111111100000000000000111110000000000000000000000000000000000000000000000000 ;
assign r_102 = 200'b00000000000000000000000111111111111100000000000000111111000000000011111111111111111110000000000001111111111111111111100111111111111100000000000000111110000000000000000000000000000000000000000000000000 ;
assign r_103 = 200'b00000000000000000001111111111111111111110000011111111100000000000000011111111111111111111111111111111111111111111001111111111111100000000000000000001111100000000000000000000000000000000000000000000000 ;
assign r_104 = 200'b00000000000000000001111111111111111111110000011111111100000000000000011111111111111111111111111111111111111111111001111111111111100000000000000000001111100000000000000000000000000000000000000000000000 ;
assign r_105 = 200'b00000000000000011111111110000000001111111111111111110000000000000000000111111111111111111111111111111101111111111111111111111100000000000000000000000111110000000000000000000000000000000000000000000000 ;
assign r_106 = 200'b00000000000000011111111110000000001111111111111111110000000000000000000111111111111111111111111111111101111111111111111111111100000000000000000000000111110000000000000000000000000000000000000000000000 ;
assign r_107 = 200'b00000000000011111111000000000000000001111111111111111110000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000011110000000000000000000000000000000000000000000000 ;
assign r_108 = 200'b00000000000011111111000000000000000001111111111111111110000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000011110000000000000000000000000000000000000000000000 ;
assign r_109 = 200'b00000000011111110000000000000000011111111111111111111111111110000000000000011111110111111111111111111111111111111111100111110000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_110 = 200'b00000000011111110000000000000000011111111111111111111111111110000000000000011111110111111111111111111111111111111111100111110000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_111 = 200'b00000001111110000000000000111111111111111000000000011111111111111111000000000011111111000000000001111111111111111011100011100000000000000000000000000001111000000000000000000000000000000000000000000000 ;
assign r_112 = 200'b00000001111110000000000000111111111111111000000000011111111111111111000000000011111111000000000001111111111111111011100011100000000000000000000000000001111000000000000000000000000000000000000000000000 ;
assign r_113 = 200'b00000011111000000000111111111111110000000000000000000000001111111111111110000000111111111111111111111011111111111011100011100000000000000000000000000001111000000000000000000000000000000000000000000000 ;
assign r_114 = 200'b00000011111000000000111111111111110000000000000000000000001111111111111110000000111111111111111111111011111111111011100011100000000000000000000000000001111000000000000000000000000000000000000000000000 ;
assign r_115 = 200'b00001111000000001111111111111111100000000000000000000000000000000111111111111100000001111111111111100111111111111111100011110000000000000000000000000000111000000000000000000000000000000000000000000000 ;
assign r_116 = 200'b00001111000000001111111111111111100000000000000000000000000000000111111111111100000001111111111111100111111111111111100011110000000000000000000000000000111000000000000000000000000000000000000000000000 ;
assign r_117 = 200'b00011110001111111111110000011111111111100000000000000000000000000000000111111111100000001111100000000000111111111110000011100000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_118 = 200'b00011110001111111111110000011111111111100000000000000000000000000000000111111111100000001111100000000000111111111110000011100000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_119 = 200'b01111111111111111000000000000000111111111111000000000000000000000000001111111111111000011110000000000000000101100011111111100000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_120 = 200'b01111111111111111000000000000000111111111111000000000000000000000000001111111111111000011110000000000000000101100011111111100000000000000000000000000001110000000000000000000000000000000000000000000000 ;
assign r_121 = 200'b11111111111100000000000000000000000000011111111110000000000000000111111111110001111110011100000000000000000111111111111111110000000000000000000000000011110000000000000000000000000000000000000000000000 ;
assign r_122 = 200'b11111111111100000000000000000000000000011111111110000000000000000111111111110001111110011100000000000000000111111111111111110000000000000000000000000011110000000000000000000000000000000000000000000000 ;
assign r_123 = 200'b11111111000000000000000000000000000000000001111111111111111111111111111100000001111111111110000000111111111111111111000001111000000000000000000000000111100000000000000000000000000000000000000000000000 ;
assign r_124 = 200'b11111111000000000000000000000000000000000001111111111111111111111111111100000001111111111110000000111111111111111111000001111000000000000000000000000111100000000000000000000000000000000000000000000000 ;
assign r_125 = 200'b11110000000000000000000000000000000000000000000001111111111111111000000000000000000111111111000001111111111100000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000 ;
assign r_126 = 200'b11110000000000000000000000000000000000000000000001111111111111111000000000000000000111111111000001111111111100000000000011111100000000000000000000001111000000000000000000000000000000000000000000000000 ;
assign r_127 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100111111110000000011111111111110000000000000000000111110000000000000000000000000000000000000000000000000 ;
assign r_128 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100111111110000000011111111111110000000000000000000111110000000000000000000000000000000000000000000000000 ;
assign r_129 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100001111100000000000000011111000000000000000000000000000000000000000000000000000 ;
assign r_130 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100001111100000000000000011111000000000000000000000000000000000000000000000000000 ;
assign r_131 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011100000111111000000000111111100000000000000000000000000000000000000000000000000000 ;
assign r_132 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111011100000111111000000000111111100000000000000000000000000000000000000000000000000000 ;
assign r_133 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000011100000010111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_134 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000011100000010111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_135 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111111111111100000011100000000000111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_136 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111111111111100000011100000000000111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_137 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_138 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_139 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_140 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_141 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_142 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_143 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_144 = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;

always@(*)begin
	case(sr)
		0   : flag = r_1  [500-col];
		1   : flag = r_2  [500-col];
		2   : flag = r_3  [500-col];
        3   : flag = r_4  [500-col];
        4   : flag = r_5  [500-col];
        5   : flag = r_6  [500-col];
        6   : flag = r_7  [500-col];
        7   : flag = r_8  [500-col];
        8   : flag = r_9  [500-col];
        9   : flag = r_10 [500-col];
        10  : flag = r_11 [500-col];
        11  : flag = r_12 [500-col];
        12  : flag = r_13 [500-col];
        13  : flag = r_14 [500-col];
        14  : flag = r_15 [500-col];
        15  : flag = r_16 [500-col];
        16  : flag = r_17 [500-col];
        17  : flag = r_18 [500-col];
        18  : flag = r_19 [500-col];
        19  : flag = r_20 [500-col];
        20  : flag = r_21 [500-col];
        21  : flag = r_22 [500-col];
        22  : flag = r_23 [500-col];
        23  : flag = r_24 [500-col];
        24  : flag = r_25 [500-col];
        25  : flag = r_26 [500-col];
        26  : flag = r_27 [500-col];
        27  : flag = r_28 [500-col];
        28  : flag = r_29 [500-col];
        29  : flag = r_30 [500-col];
        30  : flag = r_31 [500-col];
        31  : flag = r_32 [500-col];
        32  : flag = r_33 [500-col];
        33  : flag = r_34 [500-col];
        34  : flag = r_35 [500-col];
        35  : flag = r_36 [500-col];
        36  : flag = r_37 [500-col];
        37  : flag = r_38 [500-col];
        38  : flag = r_39 [500-col];
        39  : flag = r_40 [500-col];
        40  : flag = r_41 [500-col];
        41  : flag = r_42 [500-col];
        42  : flag = r_43 [500-col];
        43  : flag = r_44 [500-col];
        44  : flag = r_45 [500-col];
        45  : flag = r_46 [500-col];
        46  : flag = r_47 [500-col];
        47  : flag = r_48 [500-col];
        48  : flag = r_49 [500-col];
        49  : flag = r_50 [500-col];
        50  : flag = r_51 [500-col];
        51  : flag = r_52 [500-col];
        52  : flag = r_53 [500-col];
        53  : flag = r_54 [500-col];
        54  : flag = r_55 [500-col];
        55  : flag = r_56 [500-col];
        56  : flag = r_57 [500-col];
        57  : flag = r_58 [500-col];
        58  : flag = r_59 [500-col];
        59  : flag = r_60 [500-col];
        60  : flag = r_61 [500-col];
        61  : flag = r_62 [500-col];
        62  : flag = r_63 [500-col];
        63  : flag = r_64 [500-col];
        64  : flag = r_65 [500-col];
        65  : flag = r_66 [500-col];
        66  : flag = r_67 [500-col];
        67  : flag = r_68 [500-col];
        68  : flag = r_69 [500-col];
        69  : flag = r_70 [500-col];
        70  : flag = r_71 [500-col];
        71  : flag = r_72 [500-col];
        72  : flag = r_73 [500-col];
        73  : flag = r_74 [500-col];
        74  : flag = r_75 [500-col];
        75  : flag = r_76 [500-col];
        76  : flag = r_77 [500-col];
        77  : flag = r_78 [500-col];
        78  : flag = r_79 [500-col];
        79  : flag = r_80 [500-col];
        80  : flag = r_81 [500-col];
        81  : flag = r_82 [500-col];
        82  : flag = r_83 [500-col];
        83  : flag = r_84 [500-col];
        84  : flag = r_85 [500-col];
        85  : flag = r_86 [500-col];
        86  : flag = r_87 [500-col];
        87  : flag = r_88 [500-col];
        88  : flag = r_89 [500-col];
        89  : flag = r_90 [500-col];
        90  : flag = r_91 [500-col];
        91  : flag = r_92 [500-col];
        92  : flag = r_93 [500-col];
        93  : flag = r_94 [500-col];
        94  : flag = r_95 [500-col];
        95  : flag = r_96 [500-col];
        96  : flag = r_97 [500-col];
        97  : flag = r_98 [500-col];
        98  : flag = r_99 [500-col];
        99  : flag = r_100[500-col];
        100 : flag = r_101[500-col];
        101 : flag = r_102[500-col];
        102 : flag = r_103[500-col];
        103 : flag = r_104[500-col];
        104 : flag = r_105[500-col];
        105 : flag = r_106[500-col];
        106 : flag = r_107[500-col];
        107 : flag = r_108[500-col];
        108 : flag = r_109[500-col];
        109 : flag = r_110[500-col];
        110 : flag = r_111[500-col];
        111 : flag = r_112[500-col];
        112 : flag = r_113[500-col];
        113 : flag = r_114[500-col];
        114 : flag = r_115[500-col];
        115 : flag = r_116[500-col];
        116 : flag = r_117[500-col];
        117 : flag = r_118[500-col];
        118 : flag = r_119[500-col];
        119 : flag = r_120[500-col];
        120 : flag = r_121[500-col];
        121 : flag = r_122[500-col];
        122 : flag = r_123[500-col];
        123 : flag = r_124[500-col];
        124 : flag = r_125[500-col];
        125 : flag = r_126[500-col];
        126 : flag = r_127[500-col];
        127 : flag = r_128[500-col];
        128 : flag = r_129[500-col];
        129 : flag = r_130[500-col];
        130 : flag = r_131[500-col];
        131 : flag = r_132[500-col];
        132 : flag = r_133[500-col];
        133 : flag = r_134[500-col];
        134 : flag = r_135[500-col];
        135 : flag = r_136[500-col];
        136 : flag = r_137[500-col];
        137 : flag = r_138[500-col];
        138 : flag = r_139[500-col];
        139 : flag = r_140[500-col];
        140 : flag = r_141[500-col];
        141 : flag = r_142[500-col];
        142 : flag = r_143[500-col];
        143 : flag = r_144[500-col];
	endcase
end

always@(posedge clk)begin
	if(flag)begin
		haha <=3'b000;
	end
	else haha <= 3'b111;
end
endmodule


