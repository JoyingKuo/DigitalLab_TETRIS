`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:19:56 01/08/2017 
// Design Name: 
// Module Name:    LOSE 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LOSE(clk,row,col,lose
    );

input clk;
reg flag;
input [10:0]row,col;
output reg [2:0] lose;

wire [10:0]sr;
wire [299:0] r_1, r_2,r_3,r_4,r_5,r_6,r_7,r_8,r_9,r_10,r_11,r_12,r_13,r_14,r_15,r_16,r_17,r_18,r_19,r_20;
wire [299:0] r_21,r_22,r_23,r_24,r_25,r_26,r_27,r_28,r_29,r_30,r_31,r_32,r_33,r_34,r_35,r_36,r_37,r_38,r_39,r_40;
wire [299:0] r_41,r_42,r_43,r_44,r_45,r_46,r_47,r_48,r_49,r_50,r_51,r_52,r_53,r_54,r_55,r_56,r_57,r_58,r_59,r_60;
wire [299:0] r_61,r_62,r_63,r_64,r_65,r_66,r_67,r_68,r_69,r_70,r_71,r_72,r_73,r_74,r_75,r_76,r_77,r_78,r_79,r_80;
wire [299:0] r_81,r_82,r_83,r_84,r_85,r_86,r_87,r_88,r_89,r_90,r_91,r_92,r_93,r_94,r_95,r_96,r_97,r_98,r_99,r_100;
wire [299:0] r_101,r_102,r_103,r_104,r_105,r_106,r_107,r_108,r_109,r_110,r_111,r_112,r_113,r_114,r_115,r_116,r_117,r_118,r_119,r_120;
wire [299:0] r_121,r_122,r_123,r_124,r_125,r_126,r_127,r_128,r_129,r_130,r_131,r_132,r_133,r_134,r_135,r_136,r_137,r_138,r_139,r_140;
wire [299:0] r_141,r_142,r_143,r_144,r_145,r_146,r_147,r_148,r_149,r_150,r_151,r_152,r_153,r_154,r_155,r_156,r_157,r_158,r_159,r_160;
wire [299:0] r_161,r_162,r_163,r_164,r_165,r_166,r_167,r_168,r_169,r_170,r_171,r_172,r_173,r_174,r_175,r_176,r_177,r_178,r_179,r_180;
wire [299:0] r_181,r_182,r_183,r_184,r_185,r_186,r_187,r_188,r_189,r_190,r_191,r_192,r_193,r_194,r_195,r_196,r_197,r_198,r_199,r_200;
wire [299:0] r_201,r_202,r_203,r_204,r_205,r_206,r_207,r_208,r_209,r_210,r_211,r_212,r_213,r_214,r_215,r_216,r_217,r_218,r_219,r_220;
wire [299:0] r_221,r_222,r_223,r_224,r_225,r_226,r_227,r_228,r_229,r_230,r_231,r_232,r_233,r_234,r_235,r_236,r_237,r_238,r_239,r_240;
wire [299:0] r_241,r_242,r_243,r_244,r_245,r_246,r_247,r_248,r_249,r_250,r_251,r_252;


assign sr = row-100;

assign r_1   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_2   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_3   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_4   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_5   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_6   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_7   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_8   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_9   = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_10  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_11  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_12  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_13  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_14  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_15  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_16  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_17  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_18  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_19  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_20  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_21  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_22  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_23  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_24  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_25  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_26  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_27  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_28  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_29  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_30  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_31  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_32  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_33  = 300'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_34  = 300'b000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_35  = 300'b000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_36  = 300'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000001111111111111110000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_37  = 300'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000001111111111111110000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_38  = 300'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111000000000000000100000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_39  = 300'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_40  = 300'b000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000101111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_41  = 300'b000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000101111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_42  = 300'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000001011111111111111111111111111111111111111111111111111101000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_43  = 300'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000001011111111111111111111111111111111111111111111111111101000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_44  = 300'b000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000001011111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_45  = 300'b000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000001011111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_46  = 300'b000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000101111111111111111111111111111111111111111111111111111111111111010000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_47  = 300'b000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000101111111111111111111111111111111111111111111111111111111111111010010000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_48  = 300'b000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_49  = 300'b000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_50  = 300'b000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_51  = 300'b000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_52  = 300'b000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000001101111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_53  = 300'b000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000001101111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_54  = 300'b000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_55  = 300'b000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_56  = 300'b000000000000000000000000000000000000000000000000011111111111111111111110000000000000001000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111101010000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_57  = 300'b000000000000000000000000000000000000000000000000011111111111111111111110000000000000001000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111101010010000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_58  = 300'b000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000 ;
assign r_59  = 300'b000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000010111111111111111111111111111111111111111111111111111111111111111111111111111111111110101001000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000 ;
assign r_60  = 300'b000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_61  = 300'b000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_62  = 300'b000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000100001111111111111111111100000000000000000000000000000000000000000000000000000000000000 ;
assign r_63  = 300'b000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000 ;
assign r_64  = 300'b000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000 ;
assign r_65  = 300'b000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000 ;
assign r_66  = 300'b000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000 ;
assign r_67  = 300'b000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000 ;
assign r_68  = 300'b000000000000000000000000000000000000000000011111111111111111000000000000000000000001100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_69  = 300'b000000000000000000000000000000000000000000011111111111111111000000000000000000000001100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_70  = 300'b000000000000000000000000000000000000000001111111111111111110000000000000000000010111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_71  = 300'b000000000000000000000000000000000000000001111111111111111110000000000000000000010111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000 ;
assign r_72  = 300'b000000000000000000000000000000000000000011111111111111111000000000000001000000011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_73  = 300'b000000000000000000000000000000000000000011111111111111111000000000000000000000011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_74  = 300'b000000000000000000000000000000000000000111111111111111110000000000000000000101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_75  = 300'b000000000000000000000000000000000000000111111111111111110000000000000000000101111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_76  = 300'b000000000000000000000000000000000000000111111111111111100000000000000000010011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_77  = 300'b000000000000000000000000000000000000000111111111111111100000000000000000010011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_78  = 300'b000000000000000000000000000000000000001111111111111111000100000000000000001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000 ;
assign r_79  = 300'b000000000000000000000000000000000000001111111111111111000100000000000000001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000 ;
assign r_80  = 300'b000000000000000000000000000000000000111111111111111110000000000000000000111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111010100000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_81  = 300'b000000000000000000000000000000000000111111111111111110000000000000000000111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111010100000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_82  = 300'b000000000000000000000000000000000000111111111111111100000000000000000000111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_83  = 300'b000000000000000000000000000000000000111111111111111100000000000000000000111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_84  = 300'b000000000000000000000000000000000001111111111111111000000000000000000000111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110100000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_85  = 300'b000000000000000000000000000000000001111111111111111000000000000000000000111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111110100000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_86  = 300'b000000000000000000000000000000000011111111111111110000000000000000000000011111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111100000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_87  = 300'b000000000000000000000000000000000011111111111111110000000000000000000000011111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111100000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_88  = 300'b000000000000000000000000000000000011111111111111100000000000000000001010111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111100000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_89  = 300'b000000000000000000000000000000000011111111111111100000000000000000001010111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111100000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_90  = 300'b000000000000000000000000000000000111111111111111000000000000000000000011111111111111100011111111111111111111111111111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111110000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_91  = 300'b000000000000000000000000000000000111111111111111000000000000000000000011111111111111100011111111111111111111111111111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111110000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_92  = 300'b000000000000000000000000000000000111111111111110000000000000000000000011111111111111101011111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_93  = 300'b000000000000000000000000000000000111111111111110000000000000000000000011111111111111101011111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_94  = 300'b000000000000000000000000000000001111111111111110000000000000000000000011111111111111101011111111111111111111100000000111111111111111111111111111111111110110000000000001111111111111111111111111111011111111111000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000 ;
assign r_95  = 300'b000000000000000000000000000000001111111111111110000000000000000000000011111111111111101011111111111111111111000000000111111111111111111111111111111111110110000000000001111111111111111111111111111011111111111000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000 ;
assign r_96  = 300'b000000000000000000000000000000011111111111111100000000000000000000000011111111111110111011111111111111111011000000001001111111111111111111111111111111111100000000000000011111111111111111111111111001111111111100000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000 ;
assign r_97  = 300'b000000000000000000000000000000011111111111111100000000000000000000000011111111111110111011111111111111111011000000001001111111111111111111111111111111111100000000000000011111111111111111111111111001111111111100000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000 ;
assign r_98  = 300'b000000000000000000000000000000011111111111111000000000000000000000000001111111111110111011111111111111110110000000000111111111111111111111111111111111110000000000000100010111111111111111111111110001111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_99  = 300'b000000000000000000000000000000011111111111111000000000000000000000000001111111111110111011111111111111110110000000000111111111111111111111111111111111110000000000000100010111111111111111111111110001111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_100 = 300'b000000000000000000000000000000011111111111111000000000000000000000000001111111111110110001111111111111111000000000000011111111111111111111111111111111110000001000010000001011111111111111111111111101111111111111000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000 ;
assign r_101 = 300'b000000000000000000000000000000011111111111111000000000000000000000000001111111111110110001111111111111111000000000000011111111111111111111111111111111110000001000010000001011111111111111111111111101111111111111000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000 ;
assign r_102 = 300'b000000000000000000000000000000111111111111110000000000000000000000000011111111111111110011111111111111101010000000000011111111111111111111111111111111110011000000000000111111111111111111111111111101111111111110000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000 ;
assign r_103 = 300'b000000000000000000000000000000111111111111110000000000000000000000000011111111111111110011111111111111101010000000000011111111111111111111111111111111110011000000000000111111111111111111111111111101111111111110000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000 ;
assign r_104 = 300'b000000000000000000000000000000111111111111100000000000000000000000000011111111111111100011111111111111111000000000000000111111111111111111111111111111110100000000000000001111111111111111111111110101111111111110000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_105 = 300'b000000000000000000000000000000111111111111100000000000000000000000000011111111111111100011111111111111111000000000000000111111111111111111111111111111110100000000000000001111111111111111111111110101111111111110000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_106 = 300'b000000000000000000000000000000111111111111100000000000000000000000000001111111111111000001111111111111111100000000000111111111111111111111111111111111111100010000000010111111111111111111111111101101111111111111000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000 ;
assign r_107 = 300'b000000000000000000000000000000111111111111100000000000000000000000000001111111111111000001111111111111111100000000000111111111111111111111111111111111111100010000000010111111111111111111111111101101111111111111000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000 ;
assign r_108 = 300'b000000000000000000000000000000111111111111100000000000000000000000000001111111111111110010111111111111111100000000000111111111111111111111111111111111111110000000000101111111111111111111111111101101111111111111000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000 ;
assign r_109 = 300'b000000000000000000000000000000111111111111100000000000000000000000000001111111111111110010111111111111111100000000000111111111111111111111111111111111111110000000000101111111111111111111111111101101111111111111000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000 ;
assign r_110 = 300'b000000000000000000000000000001111111111111100000000000000000000000000011111111111111110010111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_111 = 300'b000000000000000000000000000001111111111111100000000000000000000000000011111111111111110010111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111100101111111111111000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_112 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111111110000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_113 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111111001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101111111111110000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_114 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111110000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_115 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111110000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_116 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111110000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_117 = 300'b000000000000000000000000000001111111111111000000000000000000000000000011111111111111111000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111110000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_118 = 300'b000000000000000000000000000001111111111111000000000000000000000000000010111111111111111100011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111100011111111111111010000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_119 = 300'b000000000000000000000000000001111111111111000000000000000000000000000010111111111111111100011111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111100011111111111111010000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_120 = 300'b000000000000000000000000000001111111111110000000000000000000000000000010111111111111111100011111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111000111111111111111010000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_121 = 300'b000000000000000000000000000001111111111110000000000000000000000000000010111111111111111100011111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111000111111111111111010000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_122 = 300'b000000000000000000000000000001111111111110000000000000000000000000000101111111111111111111001111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111101000111111111111111000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_123 = 300'b000000000000000000000000000001111111111110000000000000000000000000000101111111111111111111001111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111101000111111111111111000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_124 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000111111111111111110000111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111010001111111111111101000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_125 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000111111111111111110000111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111010001111111111111101000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_126 = 300'b000000000000000000000000000001111111111110000000000000000000000000000010111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111100000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_127 = 300'b000000000000000000000000000001111111111110000000000000000000000000000010111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111111111100000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_128 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_129 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000 ;
assign r_130 = 300'b000000000000000000000000000001111111111110000000000000000000000000000001001111111111111111111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111100000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_131 = 300'b000000000000000000000000000001111111111110000000000000000000000000000001001111111111111111111100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111100000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_132 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000001011111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111110100000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_133 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000001011111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111110100000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_134 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000001101111111111111111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_135 = 300'b000000000000000000000000000001111111111110000000000000000000000000000000001101111111111111111110010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000 ;
assign r_136 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000110111111111111111111000011011111111111111111111111111111111100001111111111111111111111111111111111111111111110101111111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000 ;
assign r_137 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000110111111111111111111000011011111111111111111111111111111111100001111111111111111111111111111111111111111111110101111111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000 ;
assign r_138 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000011111111111111111111111000111111111111111111111111111111110110111101111111111111111111111111111111111111101001011111111111111111010000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_139 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000011111111111111111111111000111111111111111111111111111111110110111101111111111111111111111111111111111111101001011111111111111111010000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_140 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000000101111111111111111111000011011111111111111111111111111111100000001111111111111111111111111111111111111011110111111111111111111100000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_141 = 300'b000000000000000000000000000001111111111111000000000000000000000000000000000000101111111111111111111000011011111111111111111111111111111100000001111111111111111111111111111111111111011110111111111111111111100000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_142 = 300'b000000000000000000000000000001111111111111100000000000000000000000000000000000110111111111111111111110000111111111111111111111111111100000000011101111111111111111111111111111111111100101111111111111111111000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_143 = 300'b000000000000000000000000000001111111111111100000000000000000000000000000000000110111111111111111111110000111111111111111111111111111100000000011101111111111111111111111111111111111100101111111111111111111000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000 ;
assign r_144 = 300'b000000000000000000000000000000111111111111100000000000000000000000000000000000001111111111111111111111100011011111111111111111111111100000000000111111111111111111111111111111111101101011111111111111111110000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000 ;
assign r_145 = 300'b000000000000000000000000000000111111111111100000000000000000000000000000000000001111111111111111111111100011011111111111111111111111100000000000111111111111111111111111111111111101101011111111111111111110000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000 ;
assign r_146 = 300'b000000000000000000000000000000111111111111100000000000000000000000000000000000100111111111111111111111101001011111111111111111111111110000000000010111111111111111111111111111111111000111111111111111100000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_147 = 300'b000000000000000000000000000000111111111111100000000000000000000000000000000000100011111111111111111111101001011111111111111111111111110000000000010111111111111111111111111111111111000111111111111111100000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_148 = 300'b000000000000000000000000000000111111111111110000000000000000000000000000000000000010011111111111111111111100011011111111111111111111100000000000001111111111111111111111111111111000001111111111111111001001000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_149 = 300'b000000000000000000000000000000111111111111110000000000000000000000000000000000000010011111111111111111111100011011111111111111111111100000000000001111111111111111111111111111111000001111111111111111001001000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_150 = 300'b000000000000000000000000000000111111111111110000000000000000000000000000000000001001111111111111111111111110001101111111111111111111100000000000000111111111111111111111111111111100111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_151 = 300'b000000000000000000000000000000111111111111110000000000000000000000000000000000000001111111111111111111111110001101111111111111111111100000000100000111111111111111111111111111111100111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000 ;
assign r_152 = 300'b000000000000000000000000000000011111111111111000000000000000000000000000000000000000011111111111111111111111000111111111111111111111100000000000000111111111111111111111111111111000111111111111111111000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_153 = 300'b000000000000000000000000000000011111111111111000000000000000000000000000000000000000011111111111111111111111000111111111111111111111100000000000000111111111111111111111111111111000111111111111111111000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_154 = 300'b000000000000000000000000000000011111111111111000000000000000000000000000000000000000001111111111111111111111101011111111111111111111110000000000000011111111111111111111111111101000111111111111111010000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_155 = 300'b000000000000000000000000000000011111111111111000000000000000000000000000000000000010001111111111111111111111101011111111111111111111110000000000000011111111111111111111111111101000111111111111111010000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000 ;
assign r_156 = 300'b000000000000000000000000000000001111111111111100000000000000000000000000000000000000000110111111111111111111111101111111111111111111110000000000000001111111111111111111111111011011111111111111111100000001000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000 ;
assign r_157 = 300'b000000000000000000000000000000001111111111111100000000000000000000000000000000000000000110111111111111111111111101111111111111111111110000000000000001111111111111111111111111011011111111111111111100000001000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000 ;
assign r_158 = 300'b000000000000000000000000000000001111111111111110000000000000000000000000000000000000000001111111111111111111111001111111111111111111110000000000000001111111111111111111111111100111111111111111101110000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000 ;
assign r_159 = 300'b000000000000000000000000000000001111111111111110000000000000000000000000000000000000001001111111111111111111111001111111111111111111110000000000000001111111111111111111111111100111111111111111101110000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000 ;
assign r_160 = 300'b000000000000000000000000000000000111111111111111000000000000000000000000000000001000000000111111111111111111111101011111111111111111110000000000000001011111111111111111111111100011111111111111010000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_161 = 300'b000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000111111111111111111111101011111111111111111110000001000000001011111111111111111111111100011111111111111010000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_162 = 300'b000000000000000000000000000000000111111111111111100000000000000000000000000000000000000100011111111111111111111110011111111111111111111000000000000000001111111111111111111111110111111111111111110100000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_163 = 300'b000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000011111111111111111111110011111111111111111111000000000000000001111111111111111111111110111111111111111110100000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000 ;
assign r_164 = 300'b000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000001101111111111111111111110111111111111111111100000000000000010111111111111111111111110111111111111111000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_165 = 300'b000000000000000000000000000000000011111111111111100000000000000000000000000000000000001000001101111111111111111111110111111111111111111100000000000000010111111111111111111111110111111111111111000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000 ;
assign r_166 = 300'b000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000111111111111111111111000111111111111111111100000000000000010111111111111111111110110111111111111101000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_167 = 300'b000000000000000000000000000000000001111111111111110000000000000000000000000000000000000001000111111111111111111111000111111111111111111101100000000000010111111111111111111110110111111111111101000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_168 = 300'b000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000001011111111111111111100101111111111111111111000000000000001111111111111111111110011111111111111101000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_169 = 300'b000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000001011111111111111111100101111111111111111111000000000000001111111111111111111110011111111111111101000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000 ;
assign r_170 = 300'b000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000001111111111111111111100101111111111111111110001000000001011111111111111111111110011111111111111100000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_171 = 300'b000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000001111111111111111111100101111111111111111110001000000001011111111111111111111110011111111111111100000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000 ;
assign r_172 = 300'b000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000001101111111111111111110100111111111111111111100000000000011111111111111111111111001111111111111000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000 ;
assign r_173 = 300'b000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000001101111111111111111110100111111111111111111100000000000011111111111111111111111001111111111111000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000 ;
assign r_174 = 300'b000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000010111111111111111110001111111111111111111000000000000010111111111111111111101001111111111111100000000000000000000000000000000000000011111111111111110001000000000000000000000000000000000000000000000000000 ;
assign r_175 = 300'b000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000010111111111111111110001111111111111111111000000000000010111111111111111111101001111111111111100000000000000000000000000000000000000011111111111111110001000000000000000000000000000000000000000000000000000 ;
assign r_176 = 300'b000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000010111111111111111110001011111111111111111111000000000010111111111111111111111011111111111111110100010000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_177 = 300'b000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000010111111111111111110001011111111111111111111000000000010111111111111111111111011111111111111110100010000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000 ;
assign r_178 = 300'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000010111111111111111110000011111111111111111111010000000000111111111111111111111011111111111110101000100000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_179 = 300'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000010111111111111111110000011111111111111111111010000000000111111111111111111111011111111111110101000100000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_180 = 300'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000001011111111111111111110000101111111111111111111010100000001111111111111111111001011111111111110101000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_181 = 300'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000001011111111111111111110000101111111111111111111010100000001111111111111111111001011111111111110101000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000 ;
assign r_182 = 300'b000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000001011011111111111111100000111111111111111111111110100001011111111111111111111101011111111111110101000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_183 = 300'b000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000001011011111111111111100000111111111111111111111110100001011111111111111111111101011111111111110101000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_184 = 300'b000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111111111100000000111111111111111111111111111111111111111111111110101011111111111110100000001000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_185 = 300'b000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111111111100000000111111111111111111111111111111111111111111111110101011111111111110100000001000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000 ;
assign r_186 = 300'b000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000011111111111111100000001011111111111111111111111111111111111111111111110001011111111111110100000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000 ;
assign r_187 = 300'b000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000011111111111111100000001011111111111111111111111111111111111111111111110001011111111111110100000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000 ;
assign r_188 = 300'b000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000011111111111111010000001111111111111111111111111111111111111111111111110010011111111111110001000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000 ;
assign r_189 = 300'b000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000011111111111111010000001111111111111111111111111111111111111111111111110010011111111111110001000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000 ;
assign r_190 = 300'b000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000001000111111111111111010000000010111111111111111111111111111111111111111111100010001111111111110000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_191 = 300'b000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000111111111111111010000000010111111111111111111111111111111111111111111100010001111111111110000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000 ;
assign r_192 = 300'b000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000111111111111111110000000001011111111111111111111111111111111111111010001000101111111111100000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000 ;
assign r_193 = 300'b000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000111111111111111110000110001011111111111111111111111111111111111111010001000101111111111100000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000 ;
assign r_194 = 300'b000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000111111111111111100000000001111111111111111111111111111111111111101110000100011111111111100000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_195 = 300'b000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000111111111111111100000000001111111111111111111111111111111111111101110000100011111111111100000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_196 = 300'b000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000111111111111111010000000000010111111111111111111111111111111110110000000000010111111111110000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_197 = 300'b000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000111111111111111000010000000010111111111111111111111111111111110110000000000010111111111110000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_198 = 300'b000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111101010000000000000111111111111111111111111111111011100000000000001011111111100000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_199 = 300'b000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000111111111111101010000000000000111111111111111111111111111111011100000000000001011111111100000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_200 = 300'b000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000101111111111101000000000000000001111011111111111111111110111110000000000000000101111111110000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_201 = 300'b000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000101111111111101000000000000000001111011111111111111111110111110000000000000000101111111110000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_202 = 300'b000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000101111111111100000000000000000000011111110000101100011111110000000000000000000011011110100000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_203 = 300'b000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000101111111111100000000000000000000011111110000101100011111110000000000000000000011011110100000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_204 = 300'b000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000011111111101000001000000000000000000000111111111111111000000000000000000000000000111111100000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_205 = 300'b000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000011111111101000000000000000000000000000111111111111111000000000000000000000000000111111100000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_206 = 300'b000000000000000000000000000000000000000000000000000000000011111111111111111111111100001000000000000001110110110000000000000000000000000000000000000000000000000000000000000000000000001110000000000000001111111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_207 = 300'b000000000000000000000000000000000000000000000000000000000011111111111111111111111100001000000000000001110110110000000000000000000000000000000000000000000000000000000000000000000000001110000000000000001111111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_208 = 300'b000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_209 = 300'b000000000000000000000000000000000000000000000000000000010001111111111111111111111111100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_210 = 300'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_211 = 300'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_212 = 300'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_213 = 300'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_214 = 300'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_215 = 300'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_216 = 300'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_217 = 300'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_218 = 300'b000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_219 = 300'b000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_220 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_221 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_222 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_223 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_224 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_225 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_226 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_227 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_228 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_229 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_230 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_231 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_232 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_233 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_234 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_235 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_236 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_237 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_238 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_239 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_240 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_241 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_242 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_243 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_244 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_245 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_246 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_247 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_248 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_249 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_250 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_251 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
assign r_252 = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;



always@(*)begin
	case(sr)
		0   : flag = r_1  [550-col];
		1   : flag = r_2  [550-col];
		2   : flag = r_3  [550-col];
        3   : flag = r_4  [550-col];
        4   : flag = r_5  [550-col];
        5   : flag = r_6  [550-col];
        6   : flag = r_7  [550-col];
        7   : flag = r_8  [550-col];
        8   : flag = r_9  [550-col];
        9   : flag = r_10 [550-col];
        10  : flag = r_11 [550-col];
        11  : flag = r_12 [550-col];
        12  : flag = r_13 [550-col];
        13  : flag = r_14 [550-col];
        14  : flag = r_15 [550-col];
        15  : flag = r_16 [550-col];
        16  : flag = r_17 [550-col];
        17  : flag = r_18 [550-col];
        18  : flag = r_19 [550-col];
        19  : flag = r_20 [550-col];
        20  : flag = r_21 [550-col];
        21  : flag = r_22 [550-col];
        22  : flag = r_23 [550-col];
        23  : flag = r_24 [550-col];
        24  : flag = r_25 [550-col];
        25  : flag = r_26 [550-col];
        26  : flag = r_27 [550-col];
        27  : flag = r_28 [550-col];
        28  : flag = r_29 [550-col];
        29  : flag = r_30 [550-col];
        30  : flag = r_31 [550-col];
        31  : flag = r_32 [550-col];
        32  : flag = r_33 [550-col];
        33  : flag = r_34 [550-col];
        34  : flag = r_35 [550-col];
        35  : flag = r_36 [550-col];
        36  : flag = r_37 [550-col];
        37  : flag = r_38 [550-col];
        38  : flag = r_39 [550-col];
        39  : flag = r_40 [550-col];
        40  : flag = r_41 [550-col];
        41  : flag = r_42 [550-col];
        42  : flag = r_43 [550-col];
        43  : flag = r_44 [550-col];
        44  : flag = r_45 [550-col];
        45  : flag = r_46 [550-col];
        46  : flag = r_47 [550-col];
        47  : flag = r_48 [550-col];
        48  : flag = r_49 [550-col];
        49  : flag = r_50 [550-col];
        50  : flag = r_51 [550-col];
        51  : flag = r_52 [550-col];
        52  : flag = r_53 [550-col];
        53  : flag = r_54 [550-col];
        54  : flag = r_55 [550-col];
        55  : flag = r_56 [550-col];
        56  : flag = r_57 [550-col];
        57  : flag = r_58 [550-col];
        58  : flag = r_59 [550-col];
        59  : flag = r_60 [550-col];
        60  : flag = r_61 [550-col];
        61  : flag = r_62 [550-col];
        62  : flag = r_63 [550-col];
        63  : flag = r_64 [550-col];
        64  : flag = r_65 [550-col];
        65  : flag = r_66 [550-col];
        66  : flag = r_67 [550-col];
        67  : flag = r_68 [550-col];
        68  : flag = r_69 [550-col];
        69  : flag = r_70 [550-col];
        70  : flag = r_71 [550-col];
        71  : flag = r_72 [550-col];
        72  : flag = r_73 [550-col];
        73  : flag = r_74 [550-col];
        74  : flag = r_75 [550-col];
        75  : flag = r_76 [550-col];
        76  : flag = r_77 [550-col];
        77  : flag = r_78 [550-col];
        78  : flag = r_79 [550-col];
        79  : flag = r_80 [550-col];
        80  : flag = r_81 [550-col];
        81  : flag = r_82 [550-col];
        82  : flag = r_83 [550-col];
        83  : flag = r_84 [550-col];
        84  : flag = r_85 [550-col];
        85  : flag = r_86 [550-col];
        86  : flag = r_87 [550-col];
        87  : flag = r_88 [550-col];
        88  : flag = r_89 [550-col];
        89  : flag = r_90 [550-col];
        90  : flag = r_91 [550-col];
        91  : flag = r_92 [550-col];
        92  : flag = r_93 [550-col];
        93  : flag = r_94 [550-col];
        94  : flag = r_95 [550-col];
        95  : flag = r_96 [550-col];
        96  : flag = r_97 [550-col];
        97  : flag = r_98 [550-col];
        98  : flag = r_99 [550-col];
        99  : flag = r_100[550-col];
        100 : flag = r_101[550-col];
        101 : flag = r_102[550-col];
        102 : flag = r_103[550-col];
        103 : flag = r_104[550-col];
        104 : flag = r_105[550-col];
        105 : flag = r_106[550-col];
        106 : flag = r_107[550-col];
        107 : flag = r_108[550-col];
        108 : flag = r_109[550-col];
        109 : flag = r_110[550-col];
        110 : flag = r_111[550-col];
        111 : flag = r_112[550-col];
        112 : flag = r_113[550-col];
        113 : flag = r_114[550-col];
        114 : flag = r_115[550-col];
        115 : flag = r_116[550-col];
        116 : flag = r_117[550-col];
        117 : flag = r_118[550-col];
        118 : flag = r_119[550-col];
        119 : flag = r_120[550-col];
        120 : flag = r_121[550-col];
        121 : flag = r_122[550-col];
        122 : flag = r_123[550-col];
        123 : flag = r_124[550-col];
        124 : flag = r_125[550-col];
        125 : flag = r_126[550-col];
        126 : flag = r_127[550-col];
        127 : flag = r_128[550-col];
        128 : flag = r_129[550-col];
        129 : flag = r_130[550-col];
        130 : flag = r_131[550-col];
        131 : flag = r_132[550-col];
        132 : flag = r_133[550-col];
        133 : flag = r_134[550-col];
        134 : flag = r_135[550-col];
        135 : flag = r_136[550-col];
        136 : flag = r_137[550-col];
        137 : flag = r_138[550-col];
        138 : flag = r_139[550-col];
        139 : flag = r_140[550-col];
        140 : flag = r_141[550-col];
        141 : flag = r_142[550-col];
        142 : flag = r_143[550-col];
        143 : flag = r_144[550-col];
        144 : flag = r_145[550-col];
        145 : flag = r_146[550-col];
        146 : flag = r_147[550-col];
        147 : flag = r_148[550-col];
        148 : flag = r_149[550-col];
        149 : flag = r_150[550-col];
        150 : flag = r_151[550-col];
        151 : flag = r_152[550-col];
        152 : flag = r_153[550-col];
        153 : flag = r_154[550-col];
        154 : flag = r_155[550-col];
        155 : flag = r_156[550-col];
        156 : flag = r_157[550-col];
        157 : flag = r_158[550-col];
        158 : flag = r_159[550-col];
        159 : flag = r_160[550-col];
        160 : flag = r_161[550-col];
        161 : flag = r_162[550-col];
        162 : flag = r_163[550-col];
        163 : flag = r_164[550-col];
        164 : flag = r_165[550-col];
        165 : flag = r_166[550-col];
        166 : flag = r_167[550-col];
        167 : flag = r_168[550-col];
        168 : flag = r_169[550-col];
        169 : flag = r_170[550-col];
        170 : flag = r_171[550-col];
        171 : flag = r_172[550-col];
        172 : flag = r_173[550-col];
        173 : flag = r_174[550-col];
        174 : flag = r_175[550-col];
        175 : flag = r_176[550-col];
        176 : flag = r_177[550-col];
        177 : flag = r_178[550-col];
        178 : flag = r_179[550-col];
        179 : flag = r_180[550-col];
        180 : flag = r_181[550-col];
        181 : flag = r_182[550-col];
        182 : flag = r_183[550-col];
        183 : flag = r_184[550-col];
        184 : flag = r_185[550-col];
        185 : flag = r_186[550-col];
        186 : flag = r_187[550-col];
        187 : flag = r_188[550-col];
        188 : flag = r_189[550-col];
        189 : flag = r_190[550-col];
        190 : flag = r_191[550-col];
        191 : flag = r_192[550-col];
        192 : flag = r_193[550-col];
        193 : flag = r_194[550-col];
        194 : flag = r_195[550-col];
        195 : flag = r_196[550-col];
        196 : flag = r_197[550-col];
        197 : flag = r_198[550-col];
        198 : flag = r_199[550-col];
        199 : flag = r_200[550-col];
        200 : flag = r_201[550-col];
        201 : flag = r_202[550-col];
        202 : flag = r_203[550-col];
        203 : flag = r_204[550-col];
        204 : flag = r_205[550-col];
        205 : flag = r_206[550-col];
        206 : flag = r_207[550-col];
        207 : flag = r_208[550-col];
        208 : flag = r_209[550-col];
        209 : flag = r_210[550-col];
        210 : flag = r_211[550-col];
        211 : flag = r_212[550-col];
        212 : flag = r_213[550-col];
        213 : flag = r_214[550-col];
        214 : flag = r_215[550-col];
        215 : flag = r_216[550-col];
        216 : flag = r_217[550-col];
        217 : flag = r_218[550-col];
        218 : flag = r_219[550-col];
        219 : flag = r_220[550-col];
        220 : flag = r_221[550-col];
        221 : flag = r_222[550-col];
        222 : flag = r_223[550-col];
        223 : flag = r_224[550-col];
        224 : flag = r_225[550-col];
        225 : flag = r_226[550-col];
        226 : flag = r_227[550-col];
        227 : flag = r_228[550-col];
        228 : flag = r_229[550-col];
        229 : flag = r_230[550-col];
        230 : flag = r_231[550-col];
        231 : flag = r_232[550-col];
        232 : flag = r_233[550-col];
        233 : flag = r_234[550-col];
        234 : flag = r_235[550-col];
        235 : flag = r_236[550-col];
        236 : flag = r_237[550-col];
        237 : flag = r_238[550-col];
        238 : flag = r_239[550-col];
        239 : flag = r_240[550-col];
        240 : flag = r_241[550-col];
        241 : flag = r_242[550-col];
        242 : flag = r_243[550-col];
        243 : flag = r_244[550-col];
        244 : flag = r_245[550-col];
        245 : flag = r_246[550-col];
        246 : flag = r_247[550-col];
        247 : flag = r_248[550-col];
        248 : flag = r_249[550-col];
        249 : flag = r_250[550-col];
        250 : flag = r_251[550-col];
        251 : flag = r_252[550-col];
	endcase
end

always@(posedge clk)begin
	if(flag)begin
		lose <=3'b100;
	end
	else lose <= 3'b000;
end
endmodule
