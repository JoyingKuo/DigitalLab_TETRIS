`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:26:55 01/09/2017 
// Design Name: 
// Module Name:    HA1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module HA1(clk,row,col,,haha
    );

input clk;
input sw;
reg flag;
input [10:0]row,col;
output reg [2:0] haha;

wire [10:0]sr;
wire [299:0] r_1, r_2,r_3,r_4,r_5,r_6,r_7,r_8,r_9,r_10,r_11,r_12,r_13,r_14,r_15,r_16,r_17,r_18,r_19,r_20;
wire [299:0] r_21,r_22,r_23,r_24,r_25,r_26,r_27,r_28,r_29,r_30,r_31,r_32,r_33,r_34,r_35,r_36,r_37,r_38,r_39,r_40;
wire [299:0] r_41,r_42,r_43,r_44,r_45,r_46,r_47,r_48,r_49,r_50,r_51,r_52,r_53,r_54,r_55,r_56,r_57,r_58,r_59,r_60;
wire [299:0] r_61,r_62,r_63,r_64,r_65,r_66,r_67,r_68,r_69,r_70,r_71,r_72,r_73,r_74,r_75,r_76,r_77,r_78,r_79,r_80;
wire [299:0] r_81,r_82,r_83,r_84,r_85,r_86,r_87,r_88,r_89,r_90,r_91;

assign sr = row-330;

assign r_1   = 120'b000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000;
assign r_2   = 120'b000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000;
assign r_3   = 120'b000000000000000000000000000000000000000000011111111100001111111100000011111111000000000000000000000000000000000000000000;
assign r_4   = 120'b000000000000000000000000000000000000000000011111111100001111111100000011111111000000000000000000000000000000000000000000;
assign r_5   = 120'b000000000000000000000000000000000000000111111100000001111100001111000000000111111000000000000000000000000000000000000000;
assign r_6   = 120'b000000000000000000000000000000000000000111111100000001111100001111000000000111111000000000000000000000000000000000000000;
assign r_7   = 120'b000000000000000000000000000000000000111110111111111001111000000001100000000000011110000000000000000000000000000000000000;
assign r_8   = 120'b000000000000000000000000000000000000111110111111111001111000000001100000000000011110000000000000000000000000000000000000;
assign r_9   = 120'b000000000000000000000000000000000111110011110000111111111100000000110000000000000111100000000000000000000000000000000000;
assign r_10  = 120'b000000000000000000000000000000000111110011110000111111111100000000110000000000000111100000000000000000000000000000000000;
assign r_11  = 120'b000000000000000000000000000000011110000111000000111111111100000000111111111011111101110000000000000000000000000000000000;
assign r_12  = 120'b000000000000000000000000000000011110000111000000111111111100000000111111111011111101110000000000000000000000000000000000;
assign r_13  = 120'b000000000000000000000000000001111000001100000000111111100000000000110000011111111111111000000000000000000000000000000000;
assign r_14  = 120'b000000000000000000000000000001111000001100000000111111100000000000110000011111111111111000000000000000000000000000000000;
assign r_15  = 120'b000000000000000000000000000011110000001100000000000011111000000011111111000000000011101100000000000000000000000000000000;
assign r_16  = 120'b000000000000000000000000000011110000001100000000000011111000000011111111000000000011101100000000000000000000000000000000;
assign r_17  = 120'b000000000000000000000000000111000000001100000000000111111111111111111100000000000001101110000000000000000000000000000000;
assign r_18  = 120'b000000000000000000000000000111000000001100000000000111111111111111111100000000000001101110000000000000000000000000000000;
assign r_19  = 120'b000000000000000000000000001110000001111111000000001111000011111111001111111000000001100111000000000000000000000000000000;
assign r_20  = 120'b000000000000000000000000001110000001111111000000001111000011111111001111111000000001100111000000000000000000000000000000;
assign r_21  = 120'b000000000000000000000000011100000111100011111111111110000110001111111110011100000011110011000000000000000000000000000000;
assign r_22  = 120'b000000000000000000000000011100000111100011111111111110000110001111111110011100000011110011000000000000000000000000000000;
assign r_23  = 120'b000000000000000000000000111001111111100111111111111111111100001111111111111100000111111011100000000000000000000000000000;
assign r_24  = 120'b000000000000000000000000111001111111100111111111111111111100001111111111111100000111111011100000000000000000000000000000;
assign r_25  = 120'b000000000000000000000000110011100000000000000011111100011000000111100000001111111100011101100000000000000000000000000000;
assign r_26  = 120'b000000000000000000000000110011100000000000000011111100011000000111100000001111111100011101100000000000000000000000000000;
assign r_27  = 120'b000000000000000000000001110110000000000111111111111100001100011111111111111111001100001101100000000000000000000000000000;
assign r_28  = 120'b000000000000000000000001110110000000000111111111111100001100011111111111111111001100001101100000000000000000000000000000;
assign r_29  = 120'b000000000000000000000001100110000000000000011111111101111111111110000000000000001100000111111111111000000000000000000000;
assign r_30  = 120'b000000000000000000000001100110000000000000011111111101111111111110000000000000001100000111111111111000000000000000000000;
assign r_31  = 120'b000000000000000000000001100110000000000111111110011111110000000000000000000000001100000111110000001110000000000000000000;
assign r_32  = 120'b000000000000000000000001100110000000000111111110011111110000000000000000000000001100000111110000001110000000000000000000;
assign r_33  = 120'b000000000000000000000001100111100000000000001111111000000000000000000000000000001100000111100000000111000000000000000000;
assign r_34  = 120'b000000000000000000000001100111100000000000001111111000000000000000000000000000001100000111100000000111000000000000000000;
assign r_35  = 120'b000000000000000000000001100011111100011111111100000000000000000000000000000000001100000111100000000011111111111111000000;
assign r_36  = 120'b000000000000000000000001100011111100011111111100000000000000000000000000000000001100000111100000000011111111111111000000;
assign r_37  = 120'b000000000000000000000001110011001111111110000000000000000000000000000000000000011100000111100000000011100000000111111000;
assign r_38  = 120'b000000000000000000000001110011001111111110000000000000000000000000000000000000011100000111100000000011100000000111111000;
assign r_39  = 120'b000000000000000000000000110011000011110000000000000000000000000000000000000000011000000111100000000111000000000000011110;
assign r_40  = 120'b000000000000000000000000110011000011110000000000000000000000000000000000000000011000000111100000000111000000000000011110;
assign r_41  = 120'b000000000000000000000000111011000001110000000000000000000000000000000000000000111000001111000000001111111111111111111111;
assign r_42  = 120'b000000000000000000000000111011000001110000000000000000000000000000000000000000111000001111000000001111111111111111111111;
assign r_43  = 120'b000000000000000000000000011101100000011100000000000000000000000000011111111101110000001110000000111111110000000000001111;
assign r_44  = 120'b000000000000000000000000011101100000011100000000000000000000000000011111111101110000001110000000111111110000000000001111;
assign r_45  = 120'b000000000000000000001111111111100000001110000000000000000000000011111000001111100000011111111111111001100000000000000000;
assign r_46  = 120'b000000000000000000001111111111100000001110000000000000000000000011111000001111100000011111111111111001100000000000000000;
assign r_47  = 120'b000000000000000000111111111111110000000111100000000011111111111110000000000111000000111000111111000011100000000000000000;
assign r_48  = 120'b000000000000000000111111111111110000000111100000000011111111111110000000000111000000111000111111000011100000000000000000;
assign r_49  = 120'b000000000000000001110000000011111000000001111000001110000000000000000000001110000011110001111000000111000000000000000000;
assign r_50  = 120'b000000000000000001110000000011111000000001111000001110000000000000000000001110000011110001111000000111000000000000000000;
assign r_51  = 120'b000000000000000011000000000000111100000000011110011100000000000000000000111000001111100011100000001110000000000000000000;
assign r_52  = 120'b000000000000000011000000000000111100000000011110011100000000000000000000111000001111100011100000001110000000000000000000;
assign r_53  = 120'b000000000000000011000000000000011111000000000111111000000000000000000111100000111111101111000000011100000000000000000000;
assign r_54  = 120'b000000000000000011000000000000011111000000000111111000000000000000000111100000111111101111000000011100000000000000000000;
assign r_55  = 120'b000000000000000011000000000000000111100000000000111111111100011111111110001111111111111100000001111000000000000000000000;
assign r_56  = 120'b000000000000000011000000000000000111100000000000111111111100011111111110001111111111111100000001111000000000000000000000;
assign r_57  = 120'b000000000000000001100000000000001111111100000000000001111111111111000001111111111111111000011111100000000000000000000000;
assign r_58  = 120'b000000000000000001100000000000001111111100000000000001111111111111000001111111111111111000011111100000000000000000000000;
assign r_59  = 120'b000000000000000001100000000000001111111100000000000001111111111111000001111111111111111000011111100000000000000000000000;
assign r_60  = 120'b000000000000000001100000000000001111111100000000000001111111111111000001111111111111111000011111100000000000000000000000;
assign r_61  = 120'b000000000000000001110000000000011100001111111000000000000000000001111111111111111111111111111100000000000000000000000000;
assign r_62  = 120'b000000000000000001110000000000011100001111111000000000000000000001111111111111111111111111111100000000000000000000000000;
assign r_63  = 120'b000000000000111111111100000001111000000011111111111111111111111111111011111111000000000011100000000000000000000000000000;
assign r_64  = 120'b000000000000111111111100000001111000000011111111111111111111111111111011111111000000000011100000000000000000000000000000;
assign r_65  = 120'b000000001111111000001111111111100000000000011111111111111111001111111111111100000000000000110000000000000000000000000000;
assign r_66  = 120'b000000001111111000001111111111100000000000011111111111111111001111111111111100000000000000110000000000000000000000000000;
assign r_67  = 120'b000000111100000000011111111111111111000000000111111111111111111111111111111000000000000000011000000000000000000000000000;
assign r_68  = 120'b000000111100000000011111111111111111000000000111111111111111111111111111111000000000000000011000000000000000000000000000;
assign r_69  = 120'b000011100000011111111110000000001111111111100001111111001111111111111100110000000000000000011000000000000000000000000000;
assign r_70  = 120'b000011100000011111111110000000001111111111100001111111001111111111111100110000000000000000011000000000000000000000000000;
assign r_71  = 120'b001110001111111111111100000000000000000111111111000111111110001111111100110000000000000000011000000000000000000000000000;
assign r_72  = 120'b001110001111111111111100000000000000000111111111000111111110001111111100110000000000000000011000000000000000000000000000;
assign r_73  = 120'b011111111110000000011111111000000000000000111111110011100000000011111111110000000000000000111000000000000000000000000000;
assign r_74  = 120'b011111111110000000011111111000000000000000111111110011100000000011111111110000000000000000111000000000000000000000000000;
assign r_75  = 120'b111111000000000000000000111111111111111111110000111111000001111111111110111000000000000001110000000000000000000000000000;
assign r_76  = 120'b111111000000000000000000111111111111111111110000111111000001111111111110111000000000000001110000000000000000000000000000;
assign r_77  = 120'b111111000000000000000000111111111111111111110000111111000001111111111110111000000000000001110000000000000000000000000000;
assign r_78  = 120'b110000000000000000000000000000111111111000000000001111110011111110000001111100000000000011100000000000000000000000000000;
assign r_79  = 120'b110000000000000000000000000000111111111000000000001111110011111110000001111100000000000011100000000000000000000000000000;
assign r_80  = 120'b000000000000000000000000000000000000000000000000000001111111111111111111101111000000001111000000000000000000000000000000;
assign r_81  = 120'b000000000000000000000000000000000000000000000000000001111111111111111111101111000000001111000000000000000000000000000000;
assign r_82  = 120'b000000000000000000000000000000000000000000000000000000011111111111111011000011111111111100000000000000000000000000000000;
assign r_83  = 120'b000000000000000000000000000000000000000000000000000000011111111111111011000011111111111100000000000000000000000000000000;
assign r_84  = 120'b000000000000000000000000000000000000000000000000000000011101111111000111000000011111000000000000000000000000000000000000;
assign r_85  = 120'b000000000000000000000000000000000000000000000000000000011101111111000111000000011111000000000000000000000000000000000000;
assign r_86  = 120'b000000000000000000000000000000000000000000000000000000001111000000001110000000000000000000000000000000000000000000000000;
assign r_87  = 120'b000000000000000000000000000000000000000000000000000000001111000000001110000000000000000000000000000000000000000000000000;
assign r_88  = 120'b000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000;
assign r_89  = 120'b000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000;
assign r_90  = 120'b000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000;
assign r_91  = 120'b000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000;

always@(*)begin
	case(sr)
		0   : flag = r_1  [155-col];
		1   : flag = r_2  [155-col];
		2   : flag = r_3  [155-col];
        3   : flag = r_4  [155-col];
        4   : flag = r_5  [155-col];
        5   : flag = r_6  [155-col];
        6   : flag = r_7  [155-col];
        7   : flag = r_8  [155-col];
        8   : flag = r_9  [155-col];
        9   : flag = r_10 [155-col];
        10  : flag = r_11 [155-col];
        11  : flag = r_12 [155-col];
        12  : flag = r_13 [155-col];
        13  : flag = r_14 [155-col];
        14  : flag = r_15 [155-col];
        15  : flag = r_16 [155-col];
        16  : flag = r_17 [155-col];
        17  : flag = r_18 [155-col];
        18  : flag = r_19 [155-col];
        19  : flag = r_20 [155-col];
        20  : flag = r_21 [155-col];
        21  : flag = r_22 [155-col];
        22  : flag = r_23 [155-col];
        23  : flag = r_24 [155-col];
        24  : flag = r_25 [155-col];
        25  : flag = r_26 [155-col];
        26  : flag = r_27 [155-col];
        27  : flag = r_28 [155-col];
        28  : flag = r_29 [155-col];
        29  : flag = r_30 [155-col];
        30  : flag = r_31 [155-col];
        31  : flag = r_32 [155-col];
        32  : flag = r_33 [155-col];
        33  : flag = r_34 [155-col];
        34  : flag = r_35 [155-col];
        35  : flag = r_36 [155-col];
        36  : flag = r_37 [155-col];
        37  : flag = r_38 [155-col];
        38  : flag = r_39 [155-col];
        39  : flag = r_40 [155-col];
        40  : flag = r_41 [155-col];
        41  : flag = r_42 [155-col];
        42  : flag = r_43 [155-col];
        43  : flag = r_44 [155-col];
        44  : flag = r_45 [155-col];
        45  : flag = r_46 [155-col];
        46  : flag = r_47 [155-col];
        47  : flag = r_48 [155-col];
        48  : flag = r_49 [155-col];
        49  : flag = r_50 [155-col];
        50  : flag = r_51 [155-col];
        51  : flag = r_52 [155-col];
        52  : flag = r_53 [155-col];
        53  : flag = r_54 [155-col];
        54  : flag = r_55 [155-col];
        55  : flag = r_56 [155-col];
        56  : flag = r_57 [155-col];
        57  : flag = r_58 [155-col];
        58  : flag = r_59 [155-col];
        59  : flag = r_60 [155-col];
        60  : flag = r_61 [155-col];
        61  : flag = r_62 [155-col];
        62  : flag = r_63 [155-col];
        63  : flag = r_64 [155-col];
        64  : flag = r_65 [155-col];
        65  : flag = r_66 [155-col];
        66  : flag = r_67 [155-col];
        67  : flag = r_68 [155-col];
        68  : flag = r_69 [155-col];
        69  : flag = r_70 [155-col];
        70  : flag = r_71 [155-col];
        71  : flag = r_72 [155-col];
        72  : flag = r_73 [155-col];
        73  : flag = r_74 [155-col];
        74  : flag = r_75 [155-col];
        75  : flag = r_76 [155-col];
        76  : flag = r_77 [155-col];
        77  : flag = r_78 [155-col];
        78  : flag = r_79 [155-col];
        79  : flag = r_80 [155-col];
        80  : flag = r_81 [155-col];
        81  : flag = r_82 [155-col];
        82  : flag = r_83 [155-col];
        83  : flag = r_84 [155-col];
        84  : flag = r_85 [155-col];
        85  : flag = r_86 [155-col];
        86  : flag = r_87 [155-col];
        87  : flag = r_88 [155-col];
        88  : flag = r_89 [155-col];
        89  : flag = r_90 [155-col];
        90  : flag = r_91 [155-col];
	endcase
end

always@(posedge clk)begin
	if(flag)begin
		haha <=3'b000;
	end
	else haha <= 3'b111;
end
endmodule

